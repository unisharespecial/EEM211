library verilog;
use verilog.vl_types.all;
entity aaa is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        F               : out    vl_logic
    );
end aaa;

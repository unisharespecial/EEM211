library verilog;
use verilog.vl_types.all;
entity D2_4E_MXILINX_sematik is
    port(
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        E               : in     vl_logic;
        D0              : out    vl_logic;
        D1              : out    vl_logic;
        D2              : out    vl_logic;
        D3              : out    vl_logic
    );
end D2_4E_MXILINX_sematik;

library verilog;
use verilog.vl_types.all;
entity M2_1E_MXILINX_sema3 is
    port(
        D0              : in     vl_logic;
        D1              : in     vl_logic;
        E               : in     vl_logic;
        S0              : in     vl_logic;
        O               : out    vl_logic
    );
end M2_1E_MXILINX_sema3;

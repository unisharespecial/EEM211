library verilog;
use verilog.vl_types.all;
entity TEST2 is
end TEST2;

library verilog;
use verilog.vl_types.all;
entity sema01 is
    port(
        mclk            : in     vl_logic;
        F               : out    vl_logic
    );
end sema01;

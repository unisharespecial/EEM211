library verilog;
use verilog.vl_types.all;
entity test3 is
end test3;

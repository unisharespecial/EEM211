** Profile: "SCHEMATIC1-devre2"  [ G:\Yasin\yasin2-SCHEMATIC1-devre2.sim ] 

** Creating circuit file "yasin2-SCHEMATIC1-devre2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\yasin2-SCHEMATIC1.net" 


.END

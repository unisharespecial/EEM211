library verilog;
use verilog.vl_types.all;
entity FJKC_MXILINX_sema03 is
    port(
        C               : in     vl_logic;
        CLR             : in     vl_logic;
        J               : in     vl_logic;
        K               : in     vl_logic;
        Q               : out    vl_logic
    );
end FJKC_MXILINX_sema03;

library verilog;
use verilog.vl_types.all;
entity TEST is
end TEST;

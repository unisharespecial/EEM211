library verilog;
use verilog.vl_types.all;
entity Sema2test is
end Sema2test;

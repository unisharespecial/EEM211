library verilog;
use verilog.vl_types.all;
entity M4_1E_MXILINX_sema3 is
    port(
        D0              : in     vl_logic;
        D1              : in     vl_logic;
        D2              : in     vl_logic;
        D3              : in     vl_logic;
        E               : in     vl_logic;
        S0              : in     vl_logic;
        S1              : in     vl_logic;
        O               : out    vl_logic
    );
end M4_1E_MXILINX_sema3;

** Profile: "SCHEMATIC1-devre---1"  [ G:\Yasin\yasin-SCHEMATIC1-devre---1.sim ] 

** Creating circuit file "yasin-SCHEMATIC1-devre---1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\yasin-SCHEMATIC1.net" 


.END

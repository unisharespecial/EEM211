library verilog;
use verilog.vl_types.all;
entity lab4test2 is
end lab4test2;

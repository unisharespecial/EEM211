library verilog;
use verilog.vl_types.all;
entity sss is
end sss;

library verilog;
use verilog.vl_types.all;
entity Sema1Test is
end Sema1Test;

library verilog;
use verilog.vl_types.all;
entity deny3test1 is
end deny3test1;

library verilog;
use verilog.vl_types.all;
entity sematik1 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        d               : in     vl_logic;
        F               : out    vl_logic
    );
end sematik1;

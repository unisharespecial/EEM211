library verilog;
use verilog.vl_types.all;
entity sematik1 is
    port(
        mclk            : in     vl_logic;
        F               : out    vl_logic
    );
end sematik1;

library verilog;
use verilog.vl_types.all;
entity test2 is
end test2;

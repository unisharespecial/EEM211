library verilog;
use verilog.vl_types.all;
entity lab4test is
end lab4test;
